module F1_Stage(
    input logic 
);
    logic [8:0] GHR;
    logic [31:0] PC;
    
endmodule